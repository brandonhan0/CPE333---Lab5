`timescale 1ns / 1ps
module setasscache(
    input        clk,
    input        rst,
    input [31:0] address,
    input [31:0] datain,
    input               cache_write,
    input               cache_read, 
    output logic [31:0] dataout, 
    input [1:0] MEM_SIZE, 
    input MEM_SIGN, 
    input update,
    output logic hit, 
    output logic miss, 
    output logic memory_read, 
    output logic memory_write, 
    output logic [31:0] mem_rd_addr,
    output logic [31:0] mem_wr_addr,
    input [31:0] w0, 
    input [31:0] w1, 
    input [31:0] w2, 
    input [31:0] w3, 
    output logic [31:0] ow0, 
    output logic [31:0] ow1, 
    output logic [31:0] ow2, 
    output logic [31:0] ow3,
    input [31:0] IO_IN,
    output  logic IO_WR 
);