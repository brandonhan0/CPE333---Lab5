// add modified mem file
