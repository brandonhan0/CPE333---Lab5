// guys lets make this file
